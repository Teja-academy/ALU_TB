//==================================================
// Author : Tejas-Academy
// Email  : info@tejas-academy.com
// Date   : 22-03-2025
//==================================================
 
`ifndef _ALU_REG_PREDICTOR_
`define _ALU_REG_PREDICTOR_
typedef uvm_reg_predictor#(apb_seq_item) alu_reg_predictor;
`endif
