//==================================================
// Author : Tejas-Academy
// Email  : info@tejas-academy.com
// Date   : 22-03-2025
//==================================================
//==================================================
 
`ifndef _ALU_SEQR_
`define _ALU_SEQR_
typedef uvm_sequencer#(alu_trans) alu_seqr;
`endif
